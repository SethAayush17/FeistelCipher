///////////////////////////////////////////////////////////////////////////////////////////////////
//
// Module:      proc_enable_select
// Modified:    
// Version:     1.0
// Description: This module allows you to choose between using KEY[0] to advance the processor
//              or using a 10 Hz signal generated from the 50 MHz system clock using SW[5].
//              Its inputs are the buttonpress signals generated by pressing KEY[0] and the
//              50 MHz system clock. Its output provides the processor clock to the Simple
//              Computer.
//
//              ** Note that this modules uses Verilog operators and constructs that you ** 
//              ** are NOT permittedto use in your code                                  **
//
// *****************************************
// YOU MUST NOT MODIFY ANY PART OF THIS FILE
// *****************************************
//
////////////////////////////////////////////////////////////////////////////////////////////////////

module proc_enable_select (clock, reset, manual_clock, select, clock_out);
input clock, reset, manual_clock, select;
output clock_out;
wire auto_clock;

  clockdivider divider_5Hz (clock, reset, auto_clock);
  assign clock_out = (select == 1'b0) ? manual_clock :
                     (select == 1'b1) ? auto_clock : 1'bx;

endmodule

///////////////////////////////////////////////////////////////////////////////////////////////////
//
// Module:      clockdivider
// Author:      JST/KLC
// Created:     25 October 2019
// Modified:    29 November 2021
// Version:     1.2
// Description: This module generates a 10 Hz enable signal from the 50 MHz system clock.
//              To change to 5Hz, change ALL instances of "24'd4999999" to "24'd9999999"
//
//              ** Note that this modules uses Verilog operators and constructs that you ** 
//              ** are NOT permitted to use in your code                                  **
//
//
////////////////////////////////////////////////////////////////////////////////////////////////////

module clockdivider(clock, reset, enable);
	input        clock, reset;
	output       enable;

	reg   [23:0] count;

	always@(posedge clock or posedge reset) begin
		if(reset == 1'b1)
			count <= 24'd0;
		else begin
			if(count == 24'd4999999)
				count <= 24'd0;
			else
				count <= count + 24'd1;
		end
	end
	
	assign enable = (count == 24'd4999999);
	
endmodule

